*** SPICE deck for cell T_test4{sch} from library CUDA_SPICE
*** Created on Sun Nov 25, 2018 16:50:40
*** Last revised on Sun Nov 25, 2018 16:51:25
*** Written on Sun Nov 25, 2018 16:51:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include "C:\Users\Angelinia\Documents\ESE 370\Electric\22nm_HP.pm"

.global gnd

*** TOP LEVEL CELL: T_test4{sch}
Mnmos@0 net@11 net@1 net@7 gnd N L=0.044U W=0.044U
Mnmos@1 net@7 net@1 gnd gnd N L=0.044U W=0.044U
VVDC@0 net@1 gnd DC 1V AC 0V 0
VVDC@1 net@11 gnd DC 1V AC 0V 0
.END
