*** SPICE deck for cell T_test{sch} from library CUDA_SPICE
*** Created on Fri Nov 23, 2018 13:02:25
*** Last revised on Fri Nov 23, 2018 13:06:46
*** Written on Fri Nov 23, 2018 13:07:03 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include "C:\Users\Angelinia\Documents\ESE 370\Electric\22nm_HP.pm"

.global gnd

*** TOP LEVEL CELL: T_test{sch}
Mnmos@0 net@0 net@2 gnd gnd N L=0.044U W=0.044U
Rres@0 net@0 net@5 100k
VVDC@0 net@2 gnd DC 1V AC 0V 0
VVDC@1 net@5 gnd DC 0.5V AC 0V 0
.END
