*** SPICE deck for cell Tran_T_test{sch} from library CUDA_SPICE
*** Created on Sun Dec 02, 2018 23:57:59
*** Last revised on Mon Dec 03, 2018 01:01:21
*** Written on Mon Dec 03, 2018 01:01:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include "C:\Users\Angelinia\Documents\ESE 370\Electric\22nm_HP.pm"

.global gnd vdd

*** TOP LEVEL CELL: Tran_T_test{sch}
Ccap@0 net@14 net@25 1f
Mnmos@0 net@14 net@3 gnd gnd N L=0.044U W=0.044U
Mnmos@1 net@25 net@14 gnd gnd N L=0.044U W=0.044U
Mpmos@0 vdd net@3 net@14 vdd P L=0.044U W=0.1U
Mpmos@1 vdd net@14 net@25 vdd P L=0.044U W=0.1U
VVDC@0 vdd gnd DC 1V AC 0V 0
VVPulse@0 net@3 gnd pulse (0 1V 0 0.2n 0.2n 2n 4n) DC 0V AC 0V 0
.END
