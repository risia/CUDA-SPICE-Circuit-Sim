*** SPICE deck for cell Test1{sch} from library CUDA_SPICE
*** Created on Sun Nov 18, 2018 20:03:45
*** Last revised on Sun Nov 18, 2018 20:07:25
*** Written on Sun Nov 18, 2018 20:09:44 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include "C:\Users\Angelinia\Documents\ESE 370\Electric\22nm_HP.pm"

.global gnd

*** TOP LEVEL CELL: Test1{sch}
Rres@0 net@1 net@14 1
Rres@1 net@1 net@14 1
Rres@2 gnd net@1 1
Rres@3 gnd net@3 1
Rres@4 net@3 net@1 1
II_Generi@0 net@1 gnd DC 1 AC 0
VV_Generi@0 net@14 gnd DC 1 AC 0
.END
